// ========================================================
// Instruction combinations that are valid for RISC-V
// ========================================================

`define PAT_BEQ             32'b?????????????????000?????1100011
`define PAT_BNE             32'b?????????????????001?????1100011
`define PAT_BLT             32'b?????????????????100?????1100011
`define PAT_BGE             32'b?????????????????101?????1100011
`define PAT_BLTU            32'b?????????????????110?????1100011
`define PAT_BGEU            32'b?????????????????111?????1100011
`define PAT_JALR            32'b?????????????????000?????1100111
`define PAT_JAL             32'b?????????????????????????1101111
`define PAT_LUI             32'b?????????????????????????0110111
`define PAT_AUIPC           32'b?????????????????????????0010111
`define PAT_ADDI            32'b?????????????????000?????0010011
`define PAT_SLLI            32'b000000???????????001?????0010011
`define PAT_SLTI            32'b?????????????????010?????0010011
`define PAT_SLTIU           32'b?????????????????011?????0010011
`define PAT_XORI            32'b?????????????????100?????0010011
`define PAT_SRLI            32'b000000???????????101?????0010011
`define PAT_SRAI            32'b010000???????????101?????0010011
`define PAT_ORI             32'b?????????????????110?????0010011
`define PAT_ANDI            32'b?????????????????111?????0010011
`define PAT_ADD             32'b0000000??????????000?????0110011
`define PAT_SUB             32'b0100000??????????000?????0110011
`define PAT_SLL             32'b0000000??????????001?????0110011
`define PAT_SLT             32'b0000000??????????010?????0110011
`define PAT_SLTU            32'b0000000??????????011?????0110011
`define PAT_XOR             32'b0000000??????????100?????0110011
`define PAT_SRL             32'b0000000??????????101?????0110011
`define PAT_SRA             32'b0100000??????????101?????0110011
`define PAT_OR              32'b0000000??????????110?????0110011
`define PAT_AND             32'b0000000??????????111?????0110011
`define PAT_ADDIW           32'b?????????????????000?????0011011
`define PAT_SLLIW           32'b0000000??????????001?????0011011
`define PAT_SRLIW           32'b0000000??????????101?????0011011
`define PAT_SRAIW           32'b0100000??????????101?????0011011
`define PAT_ADDW            32'b0000000??????????000?????0111011
`define PAT_SUBW            32'b0100000??????????000?????0111011
`define PAT_SLLW            32'b0000000??????????001?????0111011
`define PAT_SRLW            32'b0000000??????????101?????0111011
`define PAT_SRAW            32'b0100000??????????101?????0111011
`define PAT_LB              32'b?????????????????000?????0000011
`define PAT_LH              32'b?????????????????001?????0000011
`define PAT_LW              32'b?????????????????010?????0000011
`define PAT_LD              32'b?????????????????011?????0000011
`define PAT_LBU             32'b?????????????????100?????0000011
`define PAT_LHU             32'b?????????????????101?????0000011
`define PAT_LWU             32'b?????????????????110?????0000011
`define PAT_SB              32'b?????????????????000?????0100011
`define PAT_SH              32'b?????????????????001?????0100011
`define PAT_SW              32'b?????????????????010?????0100011
`define PAT_SD              32'b?????????????????011?????0100011
`define PAT_FENCE           32'b?????????????????000?????0001111
`define PAT_FENCE_I         32'b?????????????????001?????0001111
`define PAT_MUL             32'b0000001??????????000?????0110011
`define PAT_MULH            32'b0000001??????????001?????0110011
`define PAT_MULHSU          32'b0000001??????????010?????0110011
`define PAT_MULHU           32'b0000001??????????011?????0110011
`define PAT_DIV             32'b0000001??????????100?????0110011
`define PAT_DIVU            32'b0000001??????????101?????0110011
`define PAT_REM             32'b0000001??????????110?????0110011
`define PAT_REMU            32'b0000001??????????111?????0110011
`define PAT_MULW            32'b0000001??????????000?????0111011
`define PAT_DIVW            32'b0000001??????????100?????0111011
`define PAT_DIVUW           32'b0000001??????????101?????0111011
`define PAT_REMW            32'b0000001??????????110?????0111011
`define PAT_REMUW           32'b0000001??????????111?????0111011
`define PAT_AMOADD_W        32'b00000????????????010?????0101111
`define PAT_AMOXOR_W        32'b00100????????????010?????0101111
`define PAT_AMOOR_W         32'b01000????????????010?????0101111
`define PAT_AMOAND_W        32'b01100????????????010?????0101111
`define PAT_AMOMIN_W        32'b10000????????????010?????0101111
`define PAT_AMOMAX_W        32'b10100????????????010?????0101111
`define PAT_AMOMINU_W       32'b11000????????????010?????0101111
`define PAT_AMOMAXU_W       32'b11100????????????010?????0101111
`define PAT_AMOSWAP_W       32'b00001????????????010?????0101111
`define PAT_LR_W            32'b00010??00000?????010?????0101111
`define PAT_SC_W            32'b00011????????????010?????0101111
`define PAT_AMOADD_D        32'b00000????????????011?????0101111
`define PAT_AMOXOR_D        32'b00100????????????011?????0101111
`define PAT_AMOOR_D         32'b01000????????????011?????0101111
`define PAT_AMOAND_D        32'b01100????????????011?????0101111
`define PAT_AMOMIN_D        32'b10000????????????011?????0101111
`define PAT_AMOMAX_D        32'b10100????????????011?????0101111
`define PAT_AMOMINU_D       32'b11000????????????011?????0101111
`define PAT_AMOMAXU_D       32'b11100????????????011?????0101111
`define PAT_AMOSWAP_D       32'b00001????????????011?????0101111
`define PAT_LR_D            32'b00010??00000?????011?????0101111
`define PAT_SC_D            32'b00011????????????011?????0101111
`define PAT_ECALL           32'b00000000000000000000000001110011
`define PAT_EBREAK          32'b00000000000100000000000001110011
`define PAT_URET            32'b00000000001000000000000001110011
`define PAT_SRET            32'b00010000001000000000000001110011
`define PAT_MRET            32'b00110000001000000000000001110011
`define PAT_DRET            32'b01111011001000000000000001110011
`define PAT_SFENCE_VMA      32'b0001001??????????000000001110011
`define PAT_WFI             32'b00010000010100000000000001110011
`define PAT_CSRRW           32'b?????????????????001?????1110011
`define PAT_CSRRS           32'b?????????????????010?????1110011
`define PAT_CSRRC           32'b?????????????????011?????1110011
`define PAT_CSRRWI          32'b?????????????????101?????1110011
`define PAT_CSRRSI          32'b?????????????????110?????1110011
`define PAT_CSRRCI          32'b?????????????????111?????1110011
`define PAT_FADD_S          32'b0000000??????????????????1010011
`define PAT_FSUB_S          32'b0000100??????????????????1010011
`define PAT_FMUL_S          32'b0001000??????????????????1010011
`define PAT_FDIV_S          32'b0001100??????????????????1010011
`define PAT_FSGNJ_S         32'b0010000??????????000?????1010011
`define PAT_FSGNJN_S        32'b0010000??????????001?????1010011
`define PAT_FSGNJX_S        32'b0010000??????????010?????1010011
`define PAT_FMIN_S          32'b0010100??????????000?????1010011
`define PAT_FMAX_S          32'b0010100??????????001?????1010011
`define PAT_FSQRT_S         32'b010110000000?????????????1010011
`define PAT_FADD_D          32'b0000001??????????????????1010011
`define PAT_FSUB_D          32'b0000101??????????????????1010011
`define PAT_FMUL_D          32'b0001001??????????????????1010011
`define PAT_FDIV_D          32'b0001101??????????????????1010011
`define PAT_FSGNJ_D         32'b0010001??????????000?????1010011
`define PAT_FSGNJN_D        32'b0010001??????????001?????1010011
`define PAT_FSGNJX_D        32'b0010001??????????010?????1010011
`define PAT_FMIN_D          32'b0010101??????????000?????1010011
`define PAT_FMAX_D          32'b0010101??????????001?????1010011
`define PAT_FCVT_S_D        32'b010000000001?????????????1010011
`define PAT_FCVT_D_S        32'b010000100000?????????????1010011
`define PAT_FSQRT_D         32'b010110100000?????????????1010011
`define PAT_FADD_Q          32'b0000011??????????????????1010011
`define PAT_FSUB_Q          32'b0000111??????????????????1010011
`define PAT_FMUL_Q          32'b0001011??????????????????1010011
`define PAT_FDIV_Q          32'b0001111??????????????????1010011
`define PAT_FSGNJ_Q         32'b0010011??????????000?????1010011
`define PAT_FSGNJN_Q        32'b0010011??????????001?????1010011
`define PAT_FSGNJX_Q        32'b0010011??????????010?????1010011
`define PAT_FMIN_Q          32'b0010111??????????000?????1010011
`define PAT_FMAX_Q          32'b0010111??????????001?????1010011
`define PAT_FCVT_S_Q        32'b010000000011?????????????1010011
`define PAT_FCVT_Q_S        32'b010001100000?????????????1010011
`define PAT_FCVT_D_Q        32'b010000100011?????????????1010011
`define PAT_FCVT_Q_D        32'b010001100001?????????????1010011
`define PAT_FSQRT_Q         32'b010111100000?????????????1010011
`define PAT_FLE_S           32'b1010000??????????000?????1010011
`define PAT_FLT_S           32'b1010000??????????001?????1010011
`define PAT_FEQ_S           32'b1010000??????????010?????1010011
`define PAT_FLE_D           32'b1010001??????????000?????1010011
`define PAT_FLT_D           32'b1010001??????????001?????1010011
`define PAT_FEQ_D           32'b1010001??????????010?????1010011
`define PAT_FLE_Q           32'b1010011??????????000?????1010011
`define PAT_FLT_Q           32'b1010011??????????001?????1010011
`define PAT_FEQ_Q           32'b1010011??????????010?????1010011
`define PAT_FCVT_W_S        32'b110000000000?????????????1010011
`define PAT_FCVT_WU_S       32'b110000000001?????????????1010011
`define PAT_FCVT_L_S        32'b110000000010?????????????1010011
`define PAT_FCVT_LU_S       32'b110000000011?????????????1010011
`define PAT_FMV_X_W         32'b111000000000?????000?????1010011
`define PAT_FCLASS_S        32'b111000000000?????001?????1010011
`define PAT_FCVT_W_D        32'b110000100000?????????????1010011
`define PAT_FCVT_WU_D       32'b110000100001?????????????1010011
`define PAT_FCVT_L_D        32'b110000100010?????????????1010011
`define PAT_FCVT_LU_D       32'b110000100011?????????????1010011
`define PAT_FMV_X_D         32'b111000100000?????000?????1010011
`define PAT_FCLASS_D        32'b111000100000?????001?????1010011
`define PAT_FCVT_W_Q        32'b110001100000?????????????1010011
`define PAT_FCVT_WU_Q       32'b110001100001?????????????1010011
`define PAT_FCVT_L_Q        32'b110001100010?????????????1010011
`define PAT_FCVT_LU_Q       32'b110001100011?????????????1010011
`define PAT_FMV_X_Q         32'b111001100000?????000?????1010011
`define PAT_FCLASS_Q        32'b111001100000?????001?????1010011
`define PAT_FCVT_S_W        32'b110100000000?????????????1010011
`define PAT_FCVT_S_WU       32'b110100000001?????????????1010011
`define PAT_FCVT_S_L        32'b110100000010?????????????1010011
`define PAT_FCVT_S_LU       32'b110100000011?????????????1010011
`define PAT_FMV_W_X         32'b111100000000?????000?????1010011
`define PAT_FCVT_D_W        32'b110100100000?????????????1010011
`define PAT_FCVT_D_WU       32'b110100100001?????????????1010011
`define PAT_FCVT_D_L        32'b110100100010?????????????1010011
`define PAT_FCVT_D_LU       32'b110100100011?????????????1010011
`define PAT_FMV_D_X         32'b111100100000?????000?????1010011
`define PAT_FCVT_Q_W        32'b110101100000?????????????1010011
`define PAT_FCVT_Q_WU       32'b110101100001?????????????1010011
`define PAT_FCVT_Q_L        32'b110101100010?????????????1010011
`define PAT_FCVT_Q_LU       32'b110101100011?????????????1010011
`define PAT_FMV_Q_X         32'b111101100000?????000?????1010011
`define PAT_FLW             32'b?????????????????010?????0000111
`define PAT_FLD             32'b?????????????????011?????0000111
`define PAT_FLQ             32'b?????????????????100?????0000111
`define PAT_FSW             32'b?????????????????010?????0100111
`define PAT_FSD             32'b?????????????????011?????0100111
`define PAT_FSQ             32'b?????????????????100?????0100111
`define PAT_FMADD_S         32'b?????00??????????????????1000011
`define PAT_FMSUB_S         32'b?????00??????????????????1000111
`define PAT_FNMSUB_S        32'b?????00??????????????????1001011
`define PAT_FNMADD_S        32'b?????00??????????????????1001111
`define PAT_FMADD_D         32'b?????01??????????????????1000011
`define PAT_FMSUB_D         32'b?????01??????????????????1000111
`define PAT_FNMSUB_D        32'b?????01??????????????????1001011
`define PAT_FNMADD_D        32'b?????01??????????????????1001111
`define PAT_FMADD_Q         32'b?????11??????????????????1000011
`define PAT_FMSUB_Q         32'b?????11??????????????????1000111
`define PAT_FNMSUB_Q        32'b?????11??????????????????1001011
`define PAT_FNMADD_Q        32'b?????11??????????????????1001111
`define PAT_C_ADDI4SPN      32'b????????????????000???????????00
`define PAT_C_FLD           32'b????????????????001???????????00
`define PAT_C_LW            32'b????????????????010???????????00
`define PAT_C_FLW           32'b????????????????011???????????00
`define PAT_C_FSD           32'b????????????????101???????????00
`define PAT_C_SW            32'b????????????????110???????????00
`define PAT_C_FSW           32'b????????????????111???????????00
`define PAT_C_ADDI          32'b????????????????000???????????01
`define PAT_C_JAL           32'b????????????????001???????????01
`define PAT_C_LI            32'b????????????????010???????????01
`define PAT_C_LUI           32'b????????????????011???????????01
`define PAT_C_SRLI          32'b????????????????100?00????????01
`define PAT_C_SRAI          32'b????????????????100?01????????01
`define PAT_C_ANDI          32'b????????????????100?10????????01
`define PAT_C_SUB           32'b????????????????100011???00???01
`define PAT_C_XOR           32'b????????????????100011???01???01
`define PAT_C_OR            32'b????????????????100011???10???01
`define PAT_C_AND           32'b????????????????100011???11???01
`define PAT_C_SUBW          32'b????????????????100111???00???01
`define PAT_C_ADDW          32'b????????????????100111???01???01
`define PAT_C_J             32'b????????????????101???????????01
`define PAT_C_BEQZ          32'b????????????????110???????????01
`define PAT_C_BNEZ          32'b????????????????111???????????01
`define PAT_C_SLLI          32'b????????????????000???????????10
`define PAT_C_FLDSP         32'b????????????????001???????????10
`define PAT_C_LWSP          32'b????????????????010???????????10
`define PAT_C_FLWSP         32'b????????????????011???????????10
`define PAT_C_MV            32'b????????????????1000??????????10
`define PAT_C_ADD           32'b????????????????1001??????????10
`define PAT_C_FSDSP         32'b????????????????101???????????10
`define PAT_C_SWSP          32'b????????????????110???????????10
`define PAT_C_FSWSP         32'b????????????????111???????????10
`define PAT_C_NOP           32'b????????????????0000000000000001
`define PAT_C_ADDI16SP      32'b????????????????011?00010?????01
`define PAT_C_JR            32'b????????????????1000?????0000010
`define PAT_C_JALR          32'b????????????????1001?????0000010
`define PAT_C_EBREAK        32'b????????????????1001000000000010
`define PAT_C_LD            32'b????????????????011???????????00
`define PAT_C_SD            32'b????????????????111???????????00
`define PAT_C_ADDIW         32'b????????????????001???????????01
`define PAT_C_LDSP          32'b????????????????011???????????10
`define PAT_C_SDSP          32'b????????????????111???????????10
`define PAT_C_SLLI_RV32     32'b????????????????0000??????????10
`define PAT_C_SRLI_RV32     32'b????????????????100000????????01
`define PAT_C_SRAI_RV32     32'b????????????????100001????????01
`define PAT_CUSTOM0         32'b?????????????????000?????0001011
`define PAT_CUSTOM0_RS1     32'b?????????????????010?????0001011
`define PAT_CUSTOM0_RS1_RS2 32'b?????????????????011?????0001011
`define PAT_CUSTOM0_RD      32'b?????????????????100?????0001011
`define PAT_CUSTOM0_RD_RS1  32'b?????????????????110?????0001011
`define PAT_CUSTOM0_RD_RS1_RS2 32'b?????????????????111?????0001011
`define PAT_CUSTOM1         32'b?????????????????000?????0101011
`define PAT_CUSTOM1_RS1     32'b?????????????????010?????0101011
`define PAT_CUSTOM1_RS1_RS2 32'b?????????????????011?????0101011
`define PAT_CUSTOM1_RD      32'b?????????????????100?????0101011
`define PAT_CUSTOM1_RD_RS1  32'b?????????????????110?????0101011
`define PAT_CUSTOM1_RD_RS1_RS2 32'b?????????????????111?????0101011
`define PAT_CUSTOM2         32'b?????????????????000?????1011011
`define PAT_CUSTOM2_RS1     32'b?????????????????010?????1011011
`define PAT_CUSTOM2_RS1_RS2 32'b?????????????????011?????1011011
`define PAT_CUSTOM2_RD      32'b?????????????????100?????1011011
`define PAT_CUSTOM2_RD_RS1  32'b?????????????????110?????1011011
`define PAT_CUSTOM2_RD_RS1_RS2 32'b?????????????????111?????1011011
`define PAT_CUSTOM3         32'b?????????????????000?????1111011
`define PAT_CUSTOM3_RS1     32'b?????????????????010?????1111011
`define PAT_CUSTOM3_RS1_RS2 32'b?????????????????011?????1111011
`define PAT_CUSTOM3_RD      32'b?????????????????100?????1111011
`define PAT_CUSTOM3_RD_RS1  32'b?????????????????110?????1111011
`define PAT_CUSTOM3_RD_RS1_RS2 32'b?????????????????111?????1111011
`define PAT_SLLI_RV32       32'b0000000??????????001?????0010011
`define PAT_SRLI_RV32       32'b0000000??????????101?????0010011
`define PAT_SRAI_RV32       32'b0100000??????????101?????0010011
`define PAT_FRFLAGS         32'b00000000000100000010?????1110011
`define PAT_FSFLAGS         32'b000000000001?????001?????1110011
`define PAT_FSFLAGSI        32'b000000000001?????101?????1110011
`define PAT_FRRM            32'b00000000001000000010?????1110011
`define PAT_FSRM            32'b000000000010?????001?????1110011
`define PAT_FSRMI           32'b000000000010?????101?????1110011
`define PAT_FSCSR           32'b000000000011?????001?????1110011
`define PAT_FRCSR           32'b00000000001100000010?????1110011
`define PAT_RDCYCLE         32'b11000000000000000010?????1110011
`define PAT_RDTIME          32'b11000000000100000010?????1110011
`define PAT_RDINSTRET       32'b11000000001000000010?????1110011
`define PAT_RDCYCLEH        32'b11001000000000000010?????1110011
`define PAT_RDTIMEH         32'b11001000000100000010?????1110011
`define PAT_RDINSTRETH      32'b11001000001000000010?????1110011
`define PAT_SCALL           32'b00000000000000000000000001110011
`define PAT_SBREAK          32'b00000000000100000000000001110011
`define PAT_FMV_X_S         32'b111000000000?????000?????1010011
`define PAT_FMV_S_X         32'b111100000000?????000?????1010011
`define PAT_FENCE_TSO       32'b100000110011?????000?????0001111

